.title ECE423_HW7
.options post numdgt=8
*.inc tsmc25.net
.GLOBAL VDD!
   
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dP" PMOS 

.subckt opamp VIN1 VIN2 VOUT1 VOUT2 VCMI VCMO IREF VCM
C28 0 27  5.95071719999984E-15 M=1.0 
C29 0 7  2.35465559999998E-15 M=1.0 
C30 VDD! 27  3.9892608E-15 M=1.0 
C31 0 27  4.36848E-15 M=1.0 
C32 0 22  5.73760800000001E-15 M=1.0 
C33 0 21  2.8204416E-15 M=1.0 
C34 0 8  3.0354192E-15 M=1.0 
C35 0 7  5.9784984E-15 M=1.0 
C36 VCMO 0  3.5317584E-15 M=1.0 
C37 VOUT2 27  2.3579136E-15 M=1.0 
C38 VOUT2 0  9.05510399999995E-15 M=1.0 
C39 VDD! 0  8.63294399999997E-15 M=1.0 
C40 VOUT1 27  2.5265772E-15 M=1.0 
C41 VOUT1 0  9.40940639999997E-15 M=1.0 
C42 0 26  4.4207424E-15 M=1.0 
C43 0 25  4.4365104E-15 M=1.0 
C44 0 24  4.179564E-15 M=1.0 
C45 0 23  3.2328E-15 M=1.0 
C46 0 22  6.8572188E-15 M=1.0 
C47 0 21  5.016276E-15 M=1.0 
C48 0 8  7.5944124E-15 M=1.0 
C49 0 5  5.5873044E-15 M=1.0 
C50 0 2  2.125512E-15 M=1.0 
C51 0 VCM  3.1919868E-15 M=1.0 
C52 VOUT2 0  16.449852E-15 M=1.0 
C53 VDD! 0  28.2838464E-15 M=1.0 
C54 VOUT1 0  22.008468E-15 M=1.0 
C55 IREF 0  3.8441664E-15 M=1.0 
C56 VIN2 0  4.119768E-15 M=1.0 
C57 0 22  8.4797268E-15 M=1.0 
C58 0 21  2.035656E-15 M=1.0 
C59 0 7  2.55864E-15 M=1.0 
C60 0 3  3.3126852E-15 M=1.0 
C61 0 1  3.421488E-15 M=1.0 
C62 VOUT2 0  19.6389924E-15 M=1.0 
C63 VDD! 7  4.719312E-15 M=1.0 
C64 VDD! 0  29.9706768E-15 M=1.0 
C65 VOUT1 0  13.404396E-15 M=1.0 
C66 0 27  2.1692736E-15 M=1.0 
C67 0 5  3.4034112E-15 M=1.0 
C68 VOUT2 0  14.6701728E-15 M=1.0 
C69 VDD! 27  3.074124E-15 M=1.0 
C70 VOUT1 0  14.7142512E-15 M=1.0 
C71 VOUT1 VOUT2  5.029428E-15 M=1.0 
C72 VOUT2 21  45.5549196E-15 M=1.0 
C73 VOUT2 0  125.6035212E-15 M=1.0 
C74 VOUT1 8  45.3971196E-15 M=1.0 
C75 VOUT1 0  125.616222E-15 M=1.0 
C76 VOUT2 0  3.00084848463278E-12 M=1.0 
C77 VOUT1 0  3.00084848463278E-12 M=1.0 
C78 21 VOUT2  999.824355252255E-15 M=1.0 
C79 8 VOUT1  999.824355252255E-15 M=1.0 
M80 22 VIN2 24 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M81 24 VIN2 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M82 22 VIN2 24 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M83 24 VIN2 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M84 22 VIN2 24 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M85 24 VIN2 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M86 22 VIN2 24 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M87 24 VIN2 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M88 22 VIN2 24 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M89 22 VIN1 23 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M90 23 VIN1 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M91 22 VIN1 23 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M92 23 VIN1 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M93 22 VIN1 23 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M94 23 VIN1 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M95 22 VIN1 23 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M96 23 VIN1 22 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M97 22 VIN1 23 VDD!  TSMC25DP  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M98 22 6 6 VDD!  TSMC25DP  L=419.999992118392E-9 W=3.00000010611257E-6 
+AD=1.80000003617564E-12 AS=1.80000003617564E-12 PD=4.20000014855759E-6 
+PS=4.20000014855759E-6 M=1 
M99 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M100 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M101 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M102 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M103 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M104 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M105 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M106 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M107 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M108 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M109 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M110 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M111 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M112 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M113 IREF IREF 27 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M114 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M115 27 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M116 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M117 27 IREF IREF VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M118 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M119 VDD! 27 27 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M120 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M121 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M122 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M123 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M124 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M125 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M126 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M127 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M128 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M129 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M130 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M131 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M132 7 IREF 26 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M133 26 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M134 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M135 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M136 26 IREF 7 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M137 VDD! 27 26 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M138 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M139 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M140 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M141 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M142 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M143 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M144 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M145 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M146 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M147 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M148 21 6 24 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M149 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M150 24 6 21 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M151 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M152 25 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M153 5 IREF 25 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M154 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M155 25 IREF 5 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M156 VDD! 27 25 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M157 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M158 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M159 VOUT2 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M160 VDD! 27 VOUT2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M161 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M162 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M163 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M164 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M165 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M166 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M167 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M168 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M169 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M170 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M171 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M172 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M173 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M174 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M175 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M176 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M177 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M178 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M179 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M180 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M181 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M182 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M183 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M184 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M185 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M186 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M187 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M188 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M189 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M190 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M191 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M192 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M193 8 6 23 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M194 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M195 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M196 23 6 8 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M197 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M198 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M199 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M200 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M201 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M202 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M203 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M204 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M205 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M206 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M207 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M208 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M209 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M210 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M211 22 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M212 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M213 VDD! 27 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M214 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M215 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M216 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M217 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M218 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M219 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M220 VCMO VCMO VDD! VDD!  TSMC25DP  L=419.999992118392E-9 
+W=10.0200004453654E-6 AD=6.01199992567025E-12 AS=3.60720004213833E-12 
+PD=11.2199995783158E-6 PS=720.000002729648E-9 M=1 
M221 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M222 VDD! VCMO VCMO VDD!  TSMC25DP  L=419.999992118392E-9 
+W=10.0200004453654E-6 AD=3.60720004213833E-12 AS=3.60720004213833E-12 
+PD=720.000002729648E-9 PS=720.000002729648E-9 M=1 
M223 22 VCMI VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M224 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M225 VCMO VCMO VDD! VDD!  TSMC25DP  L=419.999992118392E-9 
+W=10.0200004453654E-6 AD=3.60720004213833E-12 AS=3.60720004213833E-12 
+PD=720.000002729648E-9 PS=720.000002729648E-9 M=1 
M226 VDD! VCMI 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M227 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M228 VDD! VCMO VCMO VDD!  TSMC25DP  L=419.999992118392E-9 
+W=10.0200004453654E-6 AD=3.60720004213833E-12 AS=6.01199992567025E-12 
+PD=720.000002729648E-9 PS=11.2199995783158E-6 M=1 
M229 22 VCMI VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M230 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M231 VDD! VCMI 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M232 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M233 22 VCMI VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M234 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M235 VDD! VCMI 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M236 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M237 22 VCMI VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M238 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M239 VDD! VCMI 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M240 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M241 22 VCMI VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M242 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M243 2 2 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M244 VDD! VCMI 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M245 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M246 VDD! 2 2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M247 22 VCMI VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M248 VOUT1 27 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M249 2 2 VDD! VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M250 VDD! VCMI 22 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M251 VDD! 27 VOUT1 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M252 VDD! 2 2 VDD!  TSMC25DP  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M253 0 5 5 0  TSMC25DN  L=419.999992118392E-9 W=1.50000005305628E-6 
+AD=900.000018087821E-15 AS=900.000018087821E-15 PD=2.70000009550131E-6 
+PS=2.70000009550131E-6 M=1 
M254 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M255 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M256 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M257 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M258 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M259 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M260 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M261 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M262 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M263 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M264 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M265 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M266 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M267 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M268 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M269 VOUT2 21 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M270 0 21 VOUT2 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M271 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M272 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M273 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M274 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M275 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M276 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M277 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M278 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M279 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M280 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M281 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M282 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M283 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M284 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M285 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M286 VOUT1 8 0 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M287 0 8 VOUT1 0  TSMC25DN  L=239.99999143598E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M288 21 5 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M289 10 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M290 10 5 21 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M291 0 7 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M292 21 5 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M293 10 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M294 10 5 21 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M295 0 7 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M296 21 5 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M297 10 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M298 10 5 21 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M299 0 7 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M300 21 5 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M301 10 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M302 10 5 21 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M303 0 7 10 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M304 9 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M305 8 5 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M306 0 7 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M307 9 5 8 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M308 8 5 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M309 9 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M310 0 7 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M311 9 5 8 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M312 9 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M313 8 5 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M314 0 7 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M315 9 5 8 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M316 9 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M317 8 5 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=3.60720004213833E-12 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M318 0 7 9 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M319 9 5 8 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M320 0 7 7 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
M321 4 5 6 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
M322 0 7 4 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
M323 3 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M324 0 7 3 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M325 3 VOUT1 VCMO 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
M326 1 7 0 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=3.60720004213833E-12 PD=11.2199995783158E-6 
+PS=720.000002729648E-9 M=1 
M327 3 VCM 2 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
M328 0 7 1 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=3.60720004213833E-12 AS=6.01199992567025E-12 PD=720.000002729648E-9 
+PS=11.2199995783158E-6 M=1 
M329 1 VCM 2 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
M330 1 VOUT2 VCMO 0  TSMC25DN  L=419.999992118392E-9 W=10.0200004453654E-6 
+AD=6.01199992567025E-12 AS=6.01199992567025E-12 PD=11.2199995783158E-6 
+PS=11.2199995783158E-6 M=1 
.ends
************************

** DEFAULT SETUP ******************************
*Xop1 vg1 vg2 out1 out2 ncm ncm IREF VCM opamp
*Cin1 vg1 0 1p
*Cin2 vg1 0 1p
*Clp1 vg1 out1 1p
*Clp2 vg2 out2 1p
***********************************************

** CMFB EVALUATION SETUP **********************
Vcmtest vt 0 DC=1.78666472 AC=1V
Xop1 vg1 vg2 out1 out2 vt cmfb_out IREF VCM opamp
Xop2 vb  vb  ot1  ot2  cmfb_out nf IREC VCM opamp
***********************************************

** DIFFERENTIAL GAIN SETUP ********************
*Xop1 vg1 vg2 out1 out2 ncm1 ncm1 IREF VCM opamp
*Xop2 vg1 vg2 ot1 ot2 ncm2 ncm2 IREF VCM opamp

*Cin1 n23 vb 1p
*Cin2 n24 vb 1p
*Rgig1 n23 vb 1g
*Rgig2 n24 vb 1g
*Clp1 n23 out1 1p
*Clp2 n24 out2 1p

*Cin3 n21 vb 1p
*Cin4 n22 vb 1p
*Rgig3 n21 vb 1g
*Rgig4 n22 vb 1g
*Clp3 n21 ot1 1p
*Clp4 n22 ot2 1p
**********************************************

** SOURCES **
Vin1 vg1 0 DC=1.25V AC=.5,180
Vin2 vg2 0 DC=1.25V AC=.5,0
VD VDD! 0 DC=2.5V
Vbb vb 0 DC=1.25V

Vvcm VCM 0 DC 1V
Iiref IREF 0 64u

** SIMULATION **
.param var=1
.temp 27
.op
*.pz V(cmfb_out) Vcmtest
*.pz V(out2) Vin1
.ac dec 10 1e3 1e9
.dc Vin1 1.249 1.251 .000001
.end
