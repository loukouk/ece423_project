.title ECE423_HW7
.options post numdgt=8
*.inc tsmc25.net
.GLOBAL VDD!
   
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dP" PMOS 

.subckt opamp VIN1 VIN2 VOUT1 VOUT2 VCMI VCMO IREF VCM
C0 VOUT1 NET67  'var*1E-12' M=1.0 
C2 VOUT1 0  'var*3E-12' M=1.0 
C3 VOUT2 0  'var*3E-12' M=1.0 
C1 VOUT2 NET79  'var*1E-12' M=1.0 
MP12 NET3 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=20 
MP10 NET3 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP3 NET22 VIN2 NET3 VDD!  TSMC25DP  L=240E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=9 
MP4 NET18 VIN1 NET3 VDD!  TSMC25DP  L=240E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=9 
MP5 NET67 NET17 NET18 VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=16 
MP6 NET79 NET17 NET22 VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=16 
MP8 NET30 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP28 NET69 IREF NET30 VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP9 NET13 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP31 VOUT2 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=34 
MP26 IREF IREF NET13 VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP16 NET17 NET17 NET3 VDD!  TSMC25DP  L=420E-9 W=3E-6 AD=1.8E-12 AS=1.8E-12 
+PD=7.2E-6 PS=7.2E-6 M=1 
MP20 NET0229 NET0229 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=4 
MP19 VCMO VCMO VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=4 
MP27 NET109 IREF NET58 VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP25 NET58 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MP30 VOUT1 NET13 VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=34 
MP7 NET3 VCMI VDD! VDD!  TSMC25DP  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=12 
MN7 NET0324 NET109 0 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MN4 VCMO VOUT2 NET0324 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=1 
MN6 NET0229 VCM NET0324 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=1 
MN0 NET67 NET69 NET71 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=8 
MN1 NET71 NET109 0 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 AS=6.012E-12 
+PD=21.24E-6 PS=21.24E-6 M=8 
MN2 NET75 NET109 0 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 AS=6.012E-12 
+PD=21.24E-6 PS=21.24E-6 M=8 
MN3 NET79 NET69 NET75 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=8 
MN20 VOUT2 NET79 0 0  TSMC25DN  L=240E-9 W=10.02E-6 AD=6.012E-12 AS=6.012E-12 
+PD=21.24E-6 PS=21.24E-6 M=17 
MN5 NET69 NET69 0 0  TSMC25DN  L=420E-9 W=1.5E-6 AD=900E-15 AS=900E-15 
+PD=4.2E-6 PS=4.2E-6 M=1 
MN18 NET17 NET69 NET95 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=1 
MN11 NET95 NET109 0 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 AS=6.012E-12 
+PD=21.24E-6 PS=21.24E-6 M=1 
MN15 NET0229 VCM NET106 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=1 
MN14 VCMO VOUT1 NET106 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=1 
MN16 NET106 NET109 0 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=2 
MN17 NET109 NET109 0 0  TSMC25DN  L=420E-9 W=10.02E-6 AD=6.012E-12 
+AS=6.012E-12 PD=21.24E-6 PS=21.24E-6 M=1 
MN19 VOUT1 NET67 0 0  TSMC25DN  L=240E-9 W=10.02E-6 AD=6.012E-12 AS=6.012E-12 
+PD=21.24E-6 PS=21.24E-6 M=17 
   
   
   
.ends
************************

** DEFAULT SETUP ******************************
*Xop1 vg1 vg2 out1 out2 ncm ncm iref1 vcm opamp
*Cin1 vg1 0 1p
*Cin2 vg1 0 1p
*Clp1 vg1 out1 1p
*Clp2 vg2 out2 1p
***********************************************

** CMFB EVALUATION SETUP **********************
*SLOW
*Vcmtest vt 0 DC=1.50227407 AC=1V
*NOMINAL
Vcmtest vt 0 DC=1.78666471 AC=1V
*FAST
*Vcmtest vt 0 DC=2.06191698 AC=1V
Xop1 vg1 vg2 out1 out2 vt cmfb_out iref1 vcm opamp
Xop2 vb  vb  ot1  ot2  cmfb_out nf iref2 vcm opamp
***********************************************

** DIFFERENTIAL GAIN SETUP ********************
*Xop1 vg1 vg2 out1 out2 ncm1 ncm1 iref1 vcm opamp
*Xop2 vg1 vg2 ot1 ot2 ncm2 ncm2 iref2 vcm opamp

*Cin1 n23 vb 1p
*Cin2 n24 vb 1p
*Rgig1 n23 vb 1g
*Rgig2 n24 vb 1g
*Clp1 n23 out1 1p
*Clp2 n24 out2 1p

*Cin3 n21 vb 1p
*Cin4 n22 vb 1p
*Rgig3 n21 vb 1g
*Rgig4 n22 vb 1g
*Clp3 n21 ot1 1p
*Clp4 n22 ot2 1p
**********************************************

** SOURCES **
Vin1 vg1 0 DC=1.25V AC=.5,180
Vin2 vg2 0 DC=1.25V AC=.5,0
*Vin vg1 vg2 DC=1V
VD VDD! 0 DC=2.5V
Vbb vb 0 DC=1.25V

vvcm vcm 0 DC 1
iiref1 iref1 0 64u M=1
iiref2 iref2 0 64u M=1

** SIMULATION **
.param var=1
.temp 27
.op
*.pz V(cmfb_out) Vcmtest
*.pz V(out2) Vin1
.ac dec 10 1e3 1e9
.dc Vin1 1.249 1.251 .000001
.end
